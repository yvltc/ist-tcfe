
* forces current values to be saved
.options savecurrents

******************************************
* input voltage source
vs 1 2 0 sin(0 180 50 0 0 90)


*Envelope detector using a full wave circuit

D1 1 3 Default
D2 2 3 Default
D3 0 1 Default
D4 0 2 Default
R1 3 0 585k
C 3 0 585u

*Voltage regulator*
R2 3 4 413.63k
D5 4 0 Default1 


.model Default D
.model Default1 D (n=19)
.op
.end

.control

*makes plots in color
set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 600e-3 400e-3


*Average
meas tran v0_REGavg AVG v(4) from=400m to=600m
meas tran v0_ENVavg AVG v(3) from=400m to=600m

*max, min v0 Regulator
meas tran v0_REGmax MAX v(4) from=400m to=600m
meas tran v0_REGmin MIN v(4) from=400m to=600m

*max, min v0 Envelope
meas tran v0_ENVmax MAX v(3) from=400m to=600m
meas tran v0_ENVmin MIN v(3) from=400m to=600m

*Envelope ripple

let v0_ENVripple = v0_ENVmax - v0_ENVmin

print v0_ENVavg v0_ENVmax v0_ENVmin v0_ENVripple

*Regulator ripple

let v0_REGripple = v0_REGmax - v0_REGmin

print v0_REGavg v0_REGmax v0_REGmin v0_REGripple

*Plots

plot v(3)
hardcopy V_ENV.eps v(3)

plot v(4)
hardcopy V_REG.eps v(4)

plot v(4)-12
hardcopy v_out-12.eps v(4)-12

let cost = ((4+19)*0.1 + 998.63 + 585)
let merit = (1/(cost * (v0_REGripple + abs(v0_REGavg-12) + 1/1000000)))
print cost merit

let VoltageDeviation = v0_REGavg-12
let VoltageRipple = v0_REGripple

echo  "op_TAB"
print VoltageDeviation VoltageRipple cost merit
echo  "op_END"

quit
.endc
