options savecurrents

.param Rin=0.1k
.param R1=100k
.param R2=40k
.param Rc=0.53k
.param Re=0.1k
.param Rout=0.16k
.param Ci=730u
.param Cb=5010u
.param Co=2950u

.csparam Rin={Rin}
.csparam R1={R1}
.csparam R2={R2}
.csparam Rc={Rc}
.csparam Re={Re}
.csparam Rout={Rout}
.csparam Ci={Ci}
.csparam Cb={Cb}
.csparam Co={Co}


* PHILIPS BJT'S
.MODEL BC557A PNP(IS=2.059E-14 ISE=2.971f ISC=1.339E-14 XTI=3 BF=227.3 BR=7.69 IKF=0.08719 IKR=0.07646 XTB=1.5 VAF=37.2 VAR=11.42 VJE=0.5912 VJC=0.1 RE=0.688 RC=0.6437 RB=1 RBM=1 IRB=1E-06 CJE=1.4E-11 CJC=1.113E-11 XCJC=0.6288 FC=0.7947 NF=1.003 NR=1.007 NE=1.316 NC=1.15 MJE=0.3572 MJC=0.3414 TF=7.046E-10 TR=1m2 ITF=0.1947 VTF=5.367 XTF=4.217 EG=1.11)
.MODEL BC547A NPN(IS=1.533E-14 ISE=7.932E-16 ISC=8.305E-14 XTI=3 BF=178.7 BR=8.628 IKF=0.1216 IKR=0.1121 XTB=1.5 VAF=69.7 VAR=44.7 VJE=0.4209 VJC=0.2 RE=0.6395 RC=0.6508 RB=1 RBM=1 IRB=1E-06 CJE=1.61E-11 CJC=4.388p XCJC=0.6193 FC=0.7762 NF=1.002 NR=1.004 NE=1.436 NC=1.207 MJE=0.3071 MJC=0.2793 TF=4.995E-10 TR=1m2 ITF=0.7021 VTF=3.523 XTF=139 EG=1.11)

Vcc vcc 0 12.0
Vin in 0 0 ac 1.0 sin(0 10m 1k)
Rin in in2 {Rin}

* input coupling capacitor
Ci in2 base {Ci}

* bias circuit
R1 vcc base {R1}
R2 base 0 {R2}

* gain stage
Q1 coll base emit BC547A
Rc vcc coll {Rc}
Re emit 0 {Re}

* bypass capacitor
Cb emit 0 {Cb}


* output stage
Q2 0 coll emit2 BC557A
Rout emit2 vcc {Rout}

* output coupling capacitor
Co emit2 out {Co}

* load
RL out 0 8

.end

.control

*makes plots in color
set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op
let vce = v(coll)-v(emit)
let vbe = v(base)-v(emit)
let vo1 = v(coll)

let vec = v(emit2)
let veb = v(emit2)-v(coll)
let vo2 = v(emit2)

echo "OPngspice_TAB"
print vbe vo1 vce veb vo2 vec
echo "OPngspice_END"

 
* time analysis
*tran 1e-5 1e-2

*plot vdb(coll)
*hardcopy vo1.eps vdb(coll)


* frequency analysis
ac dec 10 10 100MEG

plot vdb(coll)
hardcopy vo1f.eps vdb(coll)

plot vdb(out)
hardcopy vo2f.eps vdb(out)

let gain = v(out)[40]/v(in)[40]

*Maximum
let maximum = vecmax(vdb(out))-3

meas ac lcofreq WHEN vdb(out) = maximum RISE = 1
meas ac ucofreq WHEN vdb(out) = maximum CROSS = LAST

let bandwidth = ucofreq-lcofreq 

*input impedance in ohm
let Zin1 = v(in2)[40]/i(Vin)[40]/(-1)
*print all


*Cost and Merit
let cost = (Rin + R1 + R2 + Re + Rc + Rout + 8)/1000 + (Ci + Cb + Co)*10^6 + 0.1*2
let merit = abs(gain)*bandwidth/(cost*lcofreq)

echo "data_TAB"
print abs(gain) abs(Zin1) cost merit lcofreq ucofreq bandwidth
echo "data_END"

echo "values_TAB"
print Rin R1 R2 Rc Re Rout Ci Cb Co
echo "values_END"

quit
.endc

.end
