*Lowest number: 95807
*Units for the values: V, mA, kOhm, mS and uF


*Values:  R1 = 1.04921233729
*R2 = 2.01121557182
*R3 = 3.04491334831
*R4 = 4.07370420497
*R5 = 3.04829678473
*R6 = 2.08879558009
*R7 = 1.01335761883
*Vs = 5.22566789497
*C = 1.04037874222
*Kb = 7.00318569445
*Kd = 8.05999483103



* NGSPICE simulation script
* BJT amp with feedback

* forces current values to be saved
.options savecurrents

.INCLUDE data1_ng.txt
.end

.control
op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

quit
.endc
