*-----------------------------------------------------------------------------
*
* To use a subcircuit, the name must begin with 'X'.  For example:
* X1 1 2 3 4 5 uA741
*
* connections:   non-inverting input
*                |  inverting input
*                |  |  positive power supply
*                |  |  |  negative power supply
*                |  |  |  |  output
*                |  |  |  |  |
.subckt uA741    1  2  3  4  5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends



.options savecurrents

Vcc vcc 0 5.0
Vee vee 0 -5.0
Vin in 0 0 ac 1.0 sin(0 10m 1k)

C1 in non_inv 110n
C2 out 0 220n

X1 non_inv inv vcc vee amp_out uA741

R1 non_inv 0 1000
R2 amp_out out 1000
R3 amp_out inv 315k
R4 inv 0 1000


.op
.end

.control


*makes plots in color
set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0



* time analysis
tran 1e-5 1e-2

hardcopy vo1.eps v(out)

* frequency analysis
ac dec 10 10 100MEG

hardcopy vo1f.eps vdb(out)
let phase_v(out) = 180/PI*ph(v(out))
hardcopy phase.eps phase_v(out)

*central frequency
meas AC maximo MAX vdb(out) from=10 to=100MEG
meas AC fO MAX_AT vdb(out) from=10 to=100MEG

let gaindb = maximo
let gain = 10^(gaindb/20)

*low and high cut-off
let threshold = maximo-3
meas AC fL WHEN vdb(out) = threshold RISE = 1
meas AC fH WHEN vdb(out) = threshold CROSS = LAST


*input impedance in ohm
let Zin = abs(v(in)[20]/vin#branch[20]/(-1))

echo "data_TAB"
print Zin
echo "data_END"

*merit figure

let gaindev = abs(gain-100)

let freqdev = abs(fO-1000)

let cost = 13323 + (1+1+330+1) + (110+220)/1000


let merit = 1/(cost*(gaindev+freqdev+0.000001))

echo "freq_TAB"
print Fl fH fO gaindb merit cost
echo "freq_END"

quit
.endc 

