 NGSPICE simulation script
* BJT amp with feedback

* forces current values to be saved
.options savecurrents

.INCLUDE data4_ng.txt

.end
.control
op

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3


hardcopy totalresponse.ps v(6) v(1)
echo totalresponse_FIG


echo "********************************************"
echo  "Frequency response"
echo "********************************************"
AC DEC 10 0.1 1MEG

let vs = v(1)
let vc = v(6)-v(8)

hardcopy frequencyresponse.ps db(v(6)) db(vs) db(vc)
echo frequencyresponse_FIG

let phase_v(6) = 180/PI*ph(v(6))
let phase_vs = 180/PI*ph(vs)
let phase_vc = 180/PI*ph(vc)

hardcopy phase.ps phase_v(6) phase_vs phase_vc 
echo phase_FIG
 
quit
.endc
